`timescale 1ns/1ps
`include "RISCV_pkg.sv"
`include "PC_Module.sv"
`include "Instruction_Memory.sv"
`include "IF_ID_REG.sv"
`include "Control_Unit.sv"
`include "ALU_Control.sv"
`include "Imm_Block.sv"
`include "Register_File.sv"
`include "LW_Stall_Unit.sv"
`include "ID_EX_REG.sv"
`include "BEQ_J_Unit.sv"
`include "ALU_Unit.sv"
`include "Forward_Unit.sv"
`include "EX_M_REG.sv"
`include "Data_Memory.sv"
`include "M_WB_REG.sv"
`include "WB_Mux.sv"
